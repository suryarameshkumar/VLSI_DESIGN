* File: INV.pex.sp
* Created: Tue Oct  4 20:42:49 2022
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.include "INV.pex.sp.pex"
.subckt INV  GND! OUT VDD! IN
* 
* IN	IN
* VDD!	VDD!
* OUT	OUT
* GND!	GND!
XD0_noxref N_GND!_D0_noxref_pos N_VDD!_D0_noxref_neg DIODENWX  AREA=9.13886e-12
+ PERIM=1.36e-05
XMMN0 N_OUT_MMN0_d N_IN_MMN0_g N_GND!_MMN0_s N_GND!_D0_noxref_pos NFET L=7e-08
+ W=2e-06 AD=1.242e-12 AS=1.22e-12 PD=5.242e-06 PS=5.22e-06 NRD=0.0845 NRS=0.081
+ M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=6.1e-07 SB=6.21e-07 SD=0
+ PANW1=5.53e-15 PANW2=3.5e-15 PANW3=3.5e-15 PANW4=3.5e-15 PANW5=3.5e-15
+ PANW6=7e-15 PANW7=1.4e-14 PANW8=1.4e-14 PANW9=2.8e-14 PANW10=4.2e-14
XMMP0 N_OUT_MMP0_d N_IN_MMP0_g N_VDD!_MMP0_s N_VDD!_D0_noxref_neg PFET L=7e-08
+ W=4.2e-06 AD=2.4822e-12 AS=2.436e-12 PD=9.582e-06 PS=9.56e-06 NRD=0.0402381
+ NRS=0.0385714 M=1 NF=1 CNR_SWITCH=1 PCCRIT=0 PAR=1 PTWELL=1 SA=5.8e-07
+ SB=5.91e-07 SD=0 PANW1=5.95e-15 PANW2=3.5e-15 PANW3=3.5e-15 PANW4=3.5e-15
+ PANW5=3.5e-15 PANW6=1.113e-14 PANW7=2.8e-14 PANW8=6.16e-13 PANW9=5.6e-14
+ PANW10=8.4e-14
*
.include "INV.pex.sp.INV.pxi"
*
.ends
*
*
